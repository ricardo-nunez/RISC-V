----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06.03.2020 13:54:31
-- Design Name: 
-- Module Name: LATCH_D - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity LATCH_D is
    Port ( RST : in STD_LOGIC;
           EN : in STD_LOGIC;
           D : in STD_LOGIC;
           Q : out STD_LOGIC);
end LATCH_D;

architecture Behavioral of LATCH_D is
begin
    process (EN, D, RST)
    begin
RESET: 
        if (RST = '1') then 
            Q <= '0';
        elsif (EN = '1') then
            Q <= D;
        end if;       
    end process;
end Behavioral;
